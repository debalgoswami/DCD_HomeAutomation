module dcd_project();
  

     